library verilog;
use verilog.vl_types.all;
entity ALU_Testbench is
end ALU_Testbench;
